module ssdec ( 

  input logic [3:0]in, 

  input logic enable, 

  output logic [6:0]out 

); 

  

  logic [6:0] SEG7 [15:0]; 

  

  assign SEG7[4'h0] = 7'b0111111; 

  assign SEG7[4'h1] = 7'b0000110; 

  assign SEG7[4'h2] = 7'b1011011; 

  assign SEG7[4'h3] = 7'b1001111; 

  assign SEG7[4'h4] = 7'b1100110; 

  assign SEG7[4'h5] = 7'b1101101; 

  assign SEG7[4'h6] = 7'b1111101; 

  assign SEG7[4'h7] = 7'b0000111; 

  assign SEG7[4'h8] = 7'b1111111; 

  assign SEG7[4'h9] = 7'b1101111; 

  assign SEG7[4'ha] = 7'b1110111; 

  assign SEG7[4'hb] = 7'b1111100; 

  assign SEG7[4'hc] = 7'b0111001; 

  assign SEG7[4'hd] = 7'b1011110; 

  assign SEG7[4'he] = 7'b1111001; 

  assign SEG7[4'hf] = 7'b1110001; 

  

  assign out = enable == 1 ? SEG7[in]: 

        7'b0000000; 

  

endmodule 